`timescale 1ns/1ps

module and_gate(input a, input b, output out);


assign out= a && b;

endmodule
